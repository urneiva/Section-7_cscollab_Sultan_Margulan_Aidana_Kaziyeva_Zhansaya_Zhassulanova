// the width of the screen in pixels
`define LINE 799 
// the height of the screen in pixels
`define SCREEN 479

// the initial horizontal position of block in pixel
`define H_INIT 148
// the initial vertical position of block in pixel
`define V_INIT 215

`define BORDER_VLEFT 464
`define BORDER_VRIGHT 15
`define BORDER_HTOP 14
`define BORDER_HBOTTOM 798
`define BORDER_HMID_TOP 134
`define BORDER_HMID_BOTTOM 148